module video_pointer(
    input wire clk,
    input wire [4:0] x,
    input wire [4:0] y,
    input wire active,

    output reg [3:0] r,
    output reg [3:0] g,
    output reg [3:0] b,
    output reg opaque
);

    wire [15:0] pointer_r_data;
    wire [10:0] pointer_r_addr = (pointer_image * 16 * 16) + (y * 16) + x;
    wire        pointer_r_clk = clk;
    wire        pointer_r_clk_enable = 1'b1;
    wire        pointer_r_enable = 1'b1;
    wire [15:0] pointer_w_data;
    wire [10:0] pointer_w_addr;
    wire        pointer_w_clk;
    wire        pointer_w_clk_enable;
    wire        pointer_w_enable;

    wire  [1:0] pointer_color_idx = {pointer_r_data[11], pointer_r_data[13]};
    reg  [11:0] pointer_palette[2:0];
    reg   [2:0] pointer_image = 0;

    initial begin
        pointer_palette[0] = 12'h000;
        pointer_palette[1] = 12'hfff;
        pointer_palette[2] = 12'hf00;
        r = 0;
        g = 0;
        b = 0;
        opaque = 0;
    end

    always @(posedge clk) begin

        if (active) begin
            if (pointer_color_idx == 2'b0) begin
                r <= 4'd0;
                g <= 4'd0;
                b <= 4'd0;
                opaque <= 1'b0;
            end else begin
                r <= pointer_palette[pointer_color_idx-1][11:8];
                g <= pointer_palette[pointer_color_idx-1][7:4];
                b <= pointer_palette[pointer_color_idx-1][3:0];
                opaque <= 1'b1;
            end
        end else begin
            r <= 4'b0000;
            g <= 4'b0000;
            b <= 4'b0000;
            opaque <= 1'b0;
        end
    end

    SB_RAM40_4K #(
        // This initialization data is generated by sprites/spritedata.go
        // from sprite image files in that directory.
        .INIT_0(256'b0101010100000000010101010000000000000000101011110000000011110100010101010000000001010101000000000000000000001010000000001111010001010101000000000101010100000000000000000000000000000000101011010101010100000000010101010000000000000000000000000000000000001010),
        .INIT_1(256'b0101010100000000010101010000001000000000110111110000000001000000010101010000000001010101000000000000000010111111000000000100000001010101000000000101010100001111000000001111111100000000110100000101010100000000010101010000101000000000111111110000000011010000),
        .INIT_2(256'b1111111100000000111111110000000010101010000000001010101000000000111111110000000011111111001101001010101000000000101010100000000011111111000000001111111100101101101010100000110110101010000000001111111100000000111111110000101110101010010011011010101000000000),
        .INIT_3(256'b1111111100000000111111110000000010101010000000001010101000000000111111110000000011111111000000001010101000000000101010100000000011111111000000001111111100000000101010100000000010101010000000001111111100000000111111110000000010101010000000001010101000000000),
        .INIT_4(256'b0101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000),
        .INIT_5(256'b0101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000),
        .INIT_6(256'b1111111111111111111111111111111110101010101010101010101010101010111111111111111111111111111111111010101010101010101010101010101011111111111111111111111111111111101010101010101010101010101010101111111111111111111111111111111110101010101010101010101010101010),
        .INIT_7(256'b1111111111111111111111111111111110101010101010101010101010101010111111111111111111111111111111111010101010101010101010101010101011111111111111111111111111111111101010101010101010101010101010101111111111111111111111111111111110101010101010101010101010101010),
        .INIT_8(256'b0101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000),
        .INIT_9(256'b0101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000),
        .INIT_A(256'b1111111111111111111111111111111110101010101010101010101010101010111111111111111111111111111111111010101010101010101010101010101011111111111111111111111111111111101010101010101010101010101010101111111111111111111111111111111110101010101010101010101010101010),
        .INIT_B(256'b1111111111111111111111111111111110101010101010101010101010101010111111111111111111111111111111111010101010101010101010101010101011111111111111111111111111111111101010101010101010101010101010101111111111111111111111111111111110101010101010101010101010101010),
        .INIT_C(256'b0101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000),
        .INIT_D(256'b0101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000),
        .INIT_E(256'b1111111111111111111111111111111110101010101010101010101010101010111111111111111111111111111111111010101010101010101010101010101011111111111111111111111111111111101010101010101010101010101010101111111111111111111111111111111110101010101010101010101010101010),
        .INIT_F(256'b1111111111111111111111111111111110101010101010101010101010101010111111111111111111111111111111111010101010101010101010101010101011111111111111111111111111111111101010101010101010101010101010101111111111111111111111111111111110101010101010101010101010101010),
        .READ_MODE(2'd3),
        .WRITE_MODE(2'd3)
    ) pointer_ram (
        .RDATA(pointer_r_data),
        .RADDR(pointer_r_addr),
        .RCLK(pointer_r_clk),
        .RCLKE(pointer_r_clk_enable),
        .RE(pointer_r_enable) //,
        //.WDATA(pointer_w_data), 
        //.WADDR(pointer_w_addr),
        //.WCLK(pointer_w_clk),
        //.WCLKE(pointer_w_clk_enable),
        //.WE(pointer_w_enable)
    );

endmodule
