module video_pointer(
    input wire clk,
    input wire [4:0] x,
    input wire [4:0] y,
    input wire active,

    output reg [3:0] r,
    output reg [3:0] g,
    output reg [3:0] b,
    output reg opaque
);

    wire [15:0] pointer_r_data;
    wire [10:0] pointer_r_addr = (pointer_image * 16 * 16) + (y * 16) + x;
    wire        pointer_r_clk = clk;
    wire        pointer_r_clk_enable = 1'b1;
    wire        pointer_r_enable = 1'b1;
    wire [15:0] pointer_w_data;
    wire [10:0] pointer_w_addr;
    wire        pointer_w_clk;
    wire        pointer_w_clk_enable;
    wire        pointer_w_enable;

    wire  [1:0] pointer_color_idx = {pointer_r_data[11], pointer_r_data[13]};
    reg  [11:0] pointer_palette[2:0];
    reg   [2:0] pointer_image = 0;

    initial begin
        pointer_palette[0] = 12'h000;
        pointer_palette[1] = 12'hfff;
        pointer_palette[2] = 12'hf00;
        r = 0;
        g = 0;
        b = 0;
        opaque = 0;
    end

    always @(posedge clk) begin

        if (active) begin
            if (pointer_color_idx == 2'b0) begin
                r <= 4'd0;
                g <= 4'd0;
                b <= 4'd0;
                opaque <= 1'b0;
            end else begin
                r <= pointer_palette[pointer_color_idx-1][11:8];
                g <= pointer_palette[pointer_color_idx-1][7:4];
                b <= pointer_palette[pointer_color_idx-1][3:0];
                opaque <= 1'b1;
            end
        end else begin
            r <= 4'b0000;
            g <= 4'b0000;
            b <= 4'b0000;
            opaque <= 1'b0;
        end
    end

    SB_RAM40_4K #(
        // This initialization data is generated by sprites/spritedata.go
        // from sprite image files in that directory.
        .INIT_0(256'b100010001000101000100010001010001000101010110101010001000010001000100010100010001000100100010010101010001000010001000100010100010001000100000000010001000101000110001000100010100010001000100000000001000100),
        .INIT_1(256'b100010001000101000100010011010100010101010110000000000001000100010001010001000100010100010101010101100000000000010001000100010100010011101111010101010101011010001000000001000100010001010001001100110101010101010101101000100000000),
        .INIT_2(256'b1010101010101010101010101010101010001000100010001000100010001000101010101010101010101111101110101000100010001000100010001000100010101010101010101010111011111011100010001101100110001000100010001010101010101010101010101110111110011000110110011000100010001000),
        .INIT_3(256'b1010101010101010101010101010101010001000100010001000100010001000101010101010101010101010101010101000100010001000100010001000100010101010101010101010101010101010100010001000100010001000100010001010101010101010101010101010101010001000100010001000100010001000),
        .INIT_4(256'b11001100110011110011001100110000000000000000110011001100111100110011001100000000000000001100110011001111001100110011000000000000000011001100110011110011001100110000000000000000),
        .INIT_5(256'b11001100110011110011001100110000000000000000110011001100111100110011001100000000000000001100110011001111001100110011000000000000000011001100110011110011001100110000000000000000),
        .INIT_6(256'b1111111111111111111111111111111111001100110011001100110011001100111111111111111111111111111111111100110011001100110011001100110011111111111111111111111111111111110011001100110011001100110011001111111111111111111111111111111111001100110011001100110011001100),
        .INIT_7(256'b1111111111111111111111111111111111001100110011001100110011001100111111111111111111111111111111111100110011001100110011001100110011111111111111111111111111111111110011001100110011001100110011001111111111111111111111111111111111001100110011001100110011001100),
        .INIT_8(256'b11001100110011110011001100110000000000000000110011001100111100110011001100000000000000001100110011001111001100110011000000000000000011001100110011110011001100110000000000000000),
        .INIT_9(256'b11001100110011110011001100110000000000000000110011001100111100110011001100000000000000001100110011001111001100110011000000000000000011001100110011110011001100110000000000000000),
        .INIT_A(256'b1111111111111111111111111111111111001100110011001100110011001100111111111111111111111111111111111100110011001100110011001100110011111111111111111111111111111111110011001100110011001100110011001111111111111111111111111111111111001100110011001100110011001100),
        .INIT_B(256'b1111111111111111111111111111111111001100110011001100110011001100111111111111111111111111111111111100110011001100110011001100110011111111111111111111111111111111110011001100110011001100110011001111111111111111111111111111111111001100110011001100110011001100),
        .INIT_C(256'b11001100110011110011001100110000000000000000110011001100111100110011001100000000000000001100110011001111001100110011000000000000000011001100110011110011001100110000000000000000),
        .INIT_D(256'b11001100110011110011001100110000000000000000110011001100111100110011001100000000000000001100110011001111001100110011000000000000000011001100110011110011001100110000000000000000),
        .INIT_E(256'b1111111111111111111111111111111111001100110011001100110011001100111111111111111111111111111111111100110011001100110011001100110011111111111111111111111111111111110011001100110011001100110011001111111111111111111111111111111111001100110011001100110011001100),
        .INIT_F(256'b1111111111111111111111111111111111001100110011001100110011001100111111111111111111111111111111111100110011001100110011001100110011111111111111111111111111111111110011001100110011001100110011001111111111111111111111111111111111001100110011001100110011001100),
        .READ_MODE(2'd3),
        .WRITE_MODE(2'd3)
    ) pointer_ram (
        .RDATA(pointer_r_data),
        .RADDR(pointer_r_addr),
        .RCLK(pointer_r_clk),
        .RCLKE(pointer_r_clk_enable),
        .RE(pointer_r_enable) //,
        //.WDATA(pointer_w_data), 
        //.WADDR(pointer_w_addr),
        //.WCLK(pointer_w_clk),
        //.WCLKE(pointer_w_clk_enable),
        //.WE(pointer_w_enable)
    );

endmodule
