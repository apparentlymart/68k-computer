module video_pointer(
    input wire clk,
    input wire [4:0] x,
    input wire [4:0] y,
    input wire active,

    output reg [3:0] r,
    output reg [3:0] g,
    output reg [3:0] b,
    output reg opaque
);

    wire [15:0] pointer_r_data;
    reg  [10:0] pointer_r_addr = 0;
    wire        pointer_r_clk = clk;
    wire        pointer_r_clk_enable = 1'b1;
    wire        pointer_r_enable = 1'b1;
    wire [15:0] pointer_w_data;
    wire [10:0] pointer_w_addr;
    wire        pointer_w_clk;
    wire        pointer_w_clk_enable;
    wire        pointer_w_enable;

    wire  [1:0] pointer_color_idx = {pointer_r_data[11], pointer_r_data[13]};
    reg  [11:0] pointer_palette[2:0];
    reg   [2:0] pointer_image = 0;

    initial begin
        pointer_palette[0] = 12'h000;
        pointer_palette[1] = 12'hfff;
        pointer_palette[2] = 12'hf00;
        r = 0;
        g = 0;
        b = 0;
        opaque = 0;
    end

    always @(posedge clk) begin

        if (active) begin
            pointer_r_addr <= (pointer_image * 16 * 16) * (y * 16) + x;

            if (pointer_color_idx == 2'b0) begin
                r <= 4'd0;
                g <= 4'd0;
                b <= 4'd0;
                opaque <= 1'b0;
            end else begin
                r <= pointer_palette[pointer_color_idx-1][11:8];
                g <= pointer_palette[pointer_color_idx-1][7:4];
                b <= pointer_palette[pointer_color_idx-1][3:0];
                opaque <= 1'b1;
            end
        end else begin
            r <= 4'b0000;
            g <= 4'b0000;
            b <= 4'b0000;
            opaque <= 1'b0;
        end
    end

    SB_RAM40_4K #(
        // This initialization data is generated by sprites/spritedata.go
        // from sprite image files in that directory.
        .INIT_0(256'b0000000000000000000000000000000010101111101011111111010011110100000000000000000000000000000000000000101000001010111101001111010000000000000000000000000000000000000000000000000010101101101011010000000000000000000000000000000000000000000000000000101000001010),
        .INIT_1(256'b0000000000000000000000100000001011011111110111110100000001000000000000000000000000000000000000001011111110111111010000000100000000000000000000000000111100001111111111111111111111010000110100000000000000000000000010100000101011111111111111111101000011010000),
        .INIT_2(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000000000000000000000000000000000000000000000000000010110100101101000011010000110100000000000000000000000000000000000010110000101101001101010011010000000000000000),
        .INIT_3(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
        .INIT_4(256'b0000000000000000000000000000000010101111101011111111010011110100000000000000000000000000000000000000101000001010111101001111010000000000000000000000000000000000000000000000000010101101101011010000000000000000000000000000000000000000000000000000101000001010),
        .INIT_5(256'b0000000000000000000000100000001011011111110111110100000001000000000000000000000000000000000000001011111110111111010000000100000000000000000000000000111100001111111111111111111111010000110100000000000000000000000010100000101011111111111111111101000011010000),
        .INIT_6(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000000000000000000000000000000000000000000000000000010110100101101000011010000110100000000000000000000000000000000000010110000101101001101010011010000000000000000),
        .INIT_7(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
        .INIT_8(256'b0000000000000000000000000000000010101111101011111111010011110100000000000000000000000000000000000000101000001010111101001111010000000000000000000000000000000000000000000000000010101101101011010000000000000000000000000000000000000000000000000000101000001010),
        .INIT_9(256'b0000000000000000000000100000001011011111110111110100000001000000000000000000000000000000000000001011111110111111010000000100000000000000000000000000111100001111111111111111111111010000110100000000000000000000000010100000101011111111111111111101000011010000),
        .INIT_A(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000000000000000000000000000000000000000000000000000010110100101101000011010000110100000000000000000000000000000000000010110000101101001101010011010000000000000000),
        .INIT_B(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
        .INIT_C(256'b0000000000000000000000000000000010101111101011111111010011110100000000000000000000000000000000000000101000001010111101001111010000000000000000000000000000000000000000000000000010101101101011010000000000000000000000000000000000000000000000000000101000001010),
        .INIT_D(256'b0000000000000000000000100000001011011111110111110100000001000000000000000000000000000000000000001011111110111111010000000100000000000000000000000000111100001111111111111111111111010000110100000000000000000000000010100000101011111111111111111101000011010000),
        .INIT_E(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000000000000000000000000000000000000000000000000000010110100101101000011010000110100000000000000000000000000000000000010110000101101001101010011010000000000000000),
        .INIT_F(256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),
        .READ_MODE(2'd3),
        .WRITE_MODE(2'd3)
    ) pointer_ram (
        .RDATA(pointer_r_data),
        .RADDR(pointer_r_addr),
        .RCLK(pointer_r_clk),
        .RCLKE(pointer_r_clk_enable),
        .RE(pointer_r_enable) //,
        //.WDATA(pointer_w_data), 
        //.WADDR(pointer_w_addr),
        //.WCLK(pointer_w_clk),
        //.WCLKE(pointer_w_clk_enable),
        //.WE(pointer_w_enable)
    );

endmodule
